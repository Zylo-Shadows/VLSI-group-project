module Testing (
    input  wire        clk,
    input  wire        rst,  // synchronous rset
    input  wire [31:0] pc_start,
    input  wire        pc_load,
    input  wire [31:0] pc_in,
    output reg  [31:0] pc_out,
    output wire [31:0] pc_plus_4,
    output wire [31:0] pc_next
);

    always @(posedge clk) begin
        if (rst) //  rset
            pc_out <= pc_start;
        else if (pc_load)
            pc_out <= pc_in;
        else
            pc_out <= pc_out + 32'd4;
    end
 // logic 
    assign pc_plus_4 = pc_out + 32'd4;
    assign pc_next   = pc_load ? pc_in : pc_plus_4;

endmodule